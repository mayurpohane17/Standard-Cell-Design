

.include sky130nm.lib

X6 net2 A net4 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X0 net2 A VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X1 net2 A VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X2 net2 B VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X3 net2 B VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X4 Y net2 VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X5 net2 A net4 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X7 net4 B VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X8 net4 B VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X9 Y net2 VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
VDD VPWR 0 1.8
VSS VGND 0 0V

Va A VGND PULSE (0 1.8 0n 0.01n 0.01n 2ns 4ns)
Vb B VGND PULSE (0 1.8 0n 0.01n 0.01n 4ns 8ns)

C1 Y 0 0.005p



.control

foreach in_delay 0.01n 0.0230506n 0.0531329n 0.122474n 0.282311n 0.650743n 1.5n
    
    * Initiating Text Files in folder text_files
    echo "input_delay:$in_delay" >> input_delay.txt
    echo "input_delay:$in_delay" >> cell_fall.txt
    echo "input_delay:$in_delay" >> cell_rise.txt
    echo "input_delay:$in_delay" >> fall_transition.txt
    echo "input_delay:$in_delay" >> rise_transition.txt

    
    let actual_rtime = $in_delay
    
    * Changing the Va Supply Rise time as per the Input Rise Time vector
    alter @Va[pulse] = [ 0 1.8 0 $&actual_rtime $&actual_rtime 2ns 4ns ]
    
    * Input Vector - Load Cap values(index2)
    foreach out_cap 0.0005p 0.00121058p 0.002931p 0.00709641p 0.0171815p 0.0415991p 0.100718p
    
        * Changing the C1 value as per the foreach list
        alter C1 $out_cap
        
        tran 1n 20ns
        run

        * Measuring Cell Fall Time @ 50% of VDD(1.8V) 
        meas tran tinfall when v(A)=0.9 FALL=1 
        meas tran tofall when v(Y)=0.9 FALL=1
        let cfall = (tofall-tinfall)/1e-9
        echo "$&cfall" >> cell_fall.txt

        * Measuring Cell Rise Time @ 50% of VDD(1.8V) 
        meas tran tinrise when v(A)=0.9 RISE=1 
        meas tran torise when v(Y)=0.9 RISE=1
        let crise = (torise-tinrise)/1e-9
        echo "$&crise" >> cell_rise.txt

        * Measuring Fall Transion Time @ 80-20% of VDD(1.8V) 
        meas tran ft1 when v(Y)=1.44 FALL=1 
        meas tran ft2 when v(Y)=0.36 FALL=1
        let fall_tran = (ft2-ft1)/1e-9
        echo "$&fall_tran" >> fall_transition.txt
        
        * Measuring Rise Transion Time @ 20-80% of VDD(1.8V) 
        meas tran rt1 when v(Y)=1.44 RISE=1 
        meas tran rt2 when v(Y)=0.36 RISE=1
        let rise_tran = (rt1-rt2)/1e-9
        echo "$&rise_tran" >> rise_transition.txt

    end
    
    * Verification of INPUT RISE TIME
    meas tran ts1 when v(A)=1.44 RISE=1 
    meas tran ts2 when v(A)=0.36 RISE=1
    meas tran ts3 when v(A)=1.44 FALL=1 
    meas tran ts4 when v(A)=0.36 FALL=1
    let RISE_IN_SLEW = (ts1-ts2)/1e-9
    let FALL_IN_SLEW = (ts4-ts3)/1e-9
    echo "actual_rise_slew:$&RISE_IN_SLEW" >> input_delay.txt
    echo "actual_fall_slew:$&FALL_IN_SLEW" >> input_delay.txt
    

   end  
.endc
.end
