
.include sky130nm.lib

X5 net3 A net1 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X0 net3 A VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X1 net3 B VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X2 net3 C VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X4 Y net3 VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X6 net1 B net2 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X7 net2 C VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X9 Y net3 VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1


VDD VPWR 0 1.8
VSS VGND 0 0V

Va A VGND PULSE (0 1.8V 0n 0.01n 0.01n 2ns 4ns)
Vb B VGND PULSE (0 1.8V 0n 0.01n 0.01n 4ns 8ns)
Vc C VGND PULSE (0 1.8V 0n 0.01n 0.01n 8ns 16ns)

CLOAD Y 0 0.00709641p

.control

tran 1 20ns

.endc
.end  
