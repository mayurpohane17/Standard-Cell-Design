


.include sky130nm.lib

X1 C A VPWR VPWR sky130_fd_pr__pfet_01v8 l=0.15u w=0.42u
X2 C B VPWR VPWR sky130_fd_pr__pfet_01v8 l=0.15u w=0.42u

X3 C B D D sky130_fd_pr__nfet_01v8 l=0.15u w=0.42u
X4 D A VGND VGND sky130_fd_pr__nfet_01v8 l=0.15u w=0.42u

X5 X C VPWR VPWR sky130_fd_pr__pfet_01v8 l=0.15u w=0.42u
X6 X C VGND VGND sky130_fd_pr__nfet_01v8 l=0.15u w=0.42u


VDD VPWR 0 3.3V
VSS VGND 0 0V

Va A VGND PULSE (0 3.3 0n 0.1n 0.1n 2n 4n)
Vb B VGND PULSE (0 3.3 0n 0.1n 0.1n 4n 8n)

.tran 1ns 20ns

.control
run
.endc
.end
