


.include sky130nm.lib

X0 net9 A1 VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X1 net9 A2 VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X2 net9 A3 VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X3 Y B1 net9 VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X4 Y B2 net9 VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X5 Y A1 net3 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X6 net3 A2 net4 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X7 net4 A3 VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X8 Y B1 net6 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X9 net6 B2 VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1

VDD VPWR 0 1.8
VSS VGND 0 0V

Va1 A1 VGND PULSE (0 1.8 0n 0.01n 0.01n 2ns 4ns)
Va2 A2 VGND PULSE (0 1.8 0n 0.01n 0.01n 4ns 8ns)
Va3 A3 VGND PULSE (0 1.8 0n 0.01n 0.01n 8ns 16ns)
Vb1 B1 VGND PULSE (0 1.8 0n 0.01n 0.01n 16ns 32ns)
Vb2 B2 VGND PULSE (0 1.8 0n 0.01n 0.01n 32ns 64ns)

C1 Y 0 0.005p



.control

tran 1 70ns

.endc
.end
