

.include sky130nm.lib

X5 net1 A net2 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X0 net1 A VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X1 net1 B VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X2 net1 C VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X3 net1 D VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X4 Y net1 VPWR VCC sky130_fd_pr__pfet_01v8 w=0.42u l=0.15u m=1
X6 net2 B net3 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X7 net3 C net4 VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X8 net4 D VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1
X9 Y net1 VGND VSS sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u m=1

VDD VPWR 0 1.8
VSS VGND 0 0V

Va A VGND PULSE (0 1.8 0n 0.01n 0.01n 2ns 4ns)
Vb B VGND PULSE (0 1.8 0n 0.01n 0.01n 4ns 8ns)
Vc C VGND PULSE (0 1.8 0n 0.01n 0.01n 8ns 16ns)
Vd D VGND PULSE (0 1.8 0n 0.01n 0.01n 16ns 32ns)

C1 Y 0 0.005p

.control
tran 1 40ns

.endc
.end
